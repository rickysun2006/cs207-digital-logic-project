/*=============================================================================
#
# Project Name   : CS207_Project_Matrix_Calculator
# File Name      : uart_rx.sv
# Module Name    : uart_rx
# University     : SUSTech
#
# Create Date    : 2025-11-23
#
# Description    :
#     Responsible for UART input (reception).
#
# Revision History:
# -----------------------------------------------------------------------------
# Ver   |   Date     |   Author       |   Description
# -----------------------------------------------------------------------------
# v1.0  | 2025-11-23 |   [Your Name]  |   Initial creation
#
#=============================================================================*/

module uart_rx (

  );

endmodule
