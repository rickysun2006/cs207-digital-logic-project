/*=============================================================================
#
# Project Name   : CS207_Project_Matrix_Calculator
# File Name      : fpga_top.sv
# Module Name    : fpga_top
# University     : SUSTech
#
# Create Date    : 2025-11-23
#
# Description    :
#     Physical top module, responsible for clock signal input, etc.; instantiates Xilinx IP cores; handles physical button debouncing.
#
# Revision History:
# -----------------------------------------------------------------------------
# Ver   |   Date     |   Author       |   Description
# -----------------------------------------------------------------------------
# v1.0  | 2025-11-23 |   [Your Name]  |   Initial creation
#
#=============================================================================*/

module fpga_top (

  );

endmodule
