module input_image_rom (
    input wire [3:0] x, // 行地址
    input wire [3:0] y, // 列地址
    output logic [3:0] data_out // 输出
);
    // ROM 存储器定义 - 10 行×12 列 = 120 个元素
    // 使用 logic 替代 reg 以便综合器优化为组合逻辑 (如果需要)
    // 这里为了方便 ALU 调用，我们将其作为参考模型，实际 ALU 内部可能直接内嵌数据以支持并行访问
    logic [3:0] rom [0:119];

    // 初始化 ROM 内容
    initial begin
        // 第 1 行: 3 7 2 9 0 5 1 8 4 6 3 2
        rom[0] = 4'd3; rom[1] = 4'd7; rom[2] = 4'd2; rom[3] = 4'd9;
        rom[4] = 4'd0; rom[5] = 4'd5; rom[6] = 4'd1; rom[7] = 4'd8;
        rom[8] = 4'd4; rom[9] = 4'd6; rom[10] = 4'd3; rom[11] = 4'd2;

        // 第 2 行: 8 1 6 4 7 3 9 0 5 2 8 1
        rom[12] = 4'd8; rom[13] = 4'd1; rom[14] = 4'd6; rom[15] = 4'd4;
        rom[16] = 4'd7; rom[17] = 4'd3; rom[18] = 4'd9; rom[19] = 4'd0;
        rom[20] = 4'd5; rom[21] = 4'd2; rom[22] = 4'd8; rom[23] = 4'd1;

        // 第 3 行: 4 9 0 2 6 8 3 5 7 1 4 9
        rom[24] = 4'd4; rom[25] = 4'd9; rom[26] = 4'd0; rom[27] = 4'd2;
        rom[28] = 4'd6; rom[29] = 4'd8; rom[30] = 4'd3; rom[31] = 4'd5;
        rom[32] = 4'd7; rom[33] = 4'd1; rom[34] = 4'd4; rom[35] = 4'd9;

        // 第 4 行: 7 3 8 5 1 4 9 2 0 6 7 3
        rom[36] = 4'd7; rom[37] = 4'd3; rom[38] = 4'd8; rom[39] = 4'd5;
        rom[40] = 4'd1; rom[41] = 4'd4; rom[42] = 4'd9; rom[43] = 4'd2;
        rom[44] = 4'd0; rom[45] = 4'd6; rom[46] = 4'd7; rom[47] = 4'd3;

        // 第 5 行: 2 6 4 0 8 7 5 3 1 9 2 4
        rom[48] = 4'd2; rom[49] = 4'd6; rom[50] = 4'd4; rom[51] = 4'd0;
        rom[52] = 4'd8; rom[53] = 4'd7; rom[54] = 4'd5; rom[55] = 4'd3;
        rom[56] = 4'd1; rom[57] = 4'd9; rom[58] = 4'd2; rom[59] = 4'd4;

        // 第 6 行: 9 0 7 3 5 2 8 6 4 1 9 0
        rom[60] = 4'd9; rom[61] = 4'd0; rom[62] = 4'd7; rom[63] = 4'd3;
        rom[64] = 4'd5; rom[65] = 4'd2; rom[66] = 4'd8; rom[67] = 4'd6;
        rom[68] = 4'd4; rom[69] = 4'd1; rom[70] = 4'd9; rom[71] = 4'd0;

        // 第 7 行: 5 8 1 6 4 9 2 7 3 0 5 8
        rom[72] = 4'd5; rom[73] = 4'd8; rom[74] = 4'd1; rom[75] = 4'd6;
        rom[76] = 4'd4; rom[77] = 4'd9; rom[78] = 4'd2; rom[79] = 4'd7;
        rom[80] = 4'd3; rom[81] = 4'd0; rom[82] = 4'd5; rom[83] = 4'd8;

        // 第 8 行: 1 4 9 2 7 0 6 8 5 3 1 4
        rom[84] = 4'd1; rom[85] = 4'd4; rom[86] = 4'd9; rom[87] = 4'd2;
        rom[88] = 4'd7; rom[89] = 4'd0; rom[90] = 4'd6; rom[91] = 4'd8;
        rom[92] = 4'd5; rom[93] = 4'd3; rom[94] = 4'd1; rom[95] = 4'd4;

        // 第 9 行: 6 2 5 8 3 1 7 4 9 0 6 2
        rom[96] = 4'd6; rom[97] = 4'd2; rom[98] = 4'd5; rom[99] = 4'd8;
        rom[100] = 4'd3; rom[101] = 4'd1; rom[102] = 4'd7; rom[103] = 4'd4;
        rom[104] = 4'd9; rom[105] = 4'd0; rom[106] = 4'd6; rom[107] = 4'd2; // Fixed missing value

        // 第 10 行: 0 7 3 9 5 6 4 1 8 2 0 7
        rom[108] = 4'd0; rom[109] = 4'd7; rom[110] = 4'd3; rom[111] = 4'd9;
        rom[112] = 4'd5; rom[113] = 4'd6; rom[114] = 4'd4; rom[115] = 4'd1;
        rom[116] = 4'd8; rom[117] = 4'd2; rom[118] = 4'd0; rom[119] = 4'd7;
    end

    // 组合逻辑读取 (模拟 ROM)
    assign data_out = rom[x*12 + y];

endmodule
