/*=============================================================================
#
# Project Name   : CS207_Project_Matrix_Calculator
# File Name      : main_fsm.sv
# Module Name    : main_fsm
# University     : SUSTech
#
# Create Date    : 2025-11-23
#
# Description    :
#     Finite State Machine (FSM).
#
# Revision History:
# -----------------------------------------------------------------------------
# Ver   |   Date     |   Author       |   Description
# -----------------------------------------------------------------------------
# v1.0  | 2025-11-23 |   [Your Name]  |   Initial creation
#
#=============================================================================*/

module main_fsm (

  );

endmodule
